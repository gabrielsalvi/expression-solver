module operativo (variaveis ...);

    `include "components/*"


    
endmodule