module operativo ();

    `include "components/*"


    
endmodule